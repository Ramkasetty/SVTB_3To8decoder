



interface intf;
  logic enable;
  logic [2:0] In;
  logic [7:0] out;
endinterface

  

  

    





























